--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   22:30:25 03/09/2015
-- Design Name:   
-- Module Name:   C:/Users/Rodrigo/Documents/Curso_ICTP/Lab_FSM_semaforo/semaforo_tb.vhd
-- Project Name:  Lab_FSM_semaforo
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: semaforo_mod
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY semaforo_tb IS
END semaforo_tb;
 
ARCHITECTURE behavior OF semaforo_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT semaforo_mod
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         red : OUT  std_logic;
         yellow : OUT  std_logic;
         green : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';

 	--Outputs
   signal red : std_logic;
   signal yellow : std_logic;
   signal green : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: semaforo_mod PORT MAP (
          clk => clk,
          rst => rst,
          red => red,
          yellow => yellow,
          green => green
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		rst <= '1';
      wait for clk_period*3;		

		rst <= '0';
      wait for clk_period*20;

      wait;
   end process;

END;
